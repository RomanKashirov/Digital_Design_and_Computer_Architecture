module mem(input  logic clk, we,
           input  logic [31:0] a, wd,
           output logic [31:0] rd);
  logic [31:0] RAM[63:0];
  initial
    $readmemh("D:/Git/Digital_Design_and_Computer_Architecture/ARM Edition/MULTICYCLE_ARM_PROCESSOR/memfile.dat",RAM);
    assign rd = RAM[a[31:2]]; // выровнять на границу слова
    always_ff @(posedge clk)
      if (we) RAM[a[31:2]] <= wd;
endmodule
