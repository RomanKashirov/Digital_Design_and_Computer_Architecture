module maindecfsm(input logic clk, reset,
						input  logic [5:0] op,
						output logic memwrite,
						output logic lord, irwrite, regdst, memtoreg,
                  output  logic regwrite, alusrca,
                  output logic [1:0]  alusrcb,
						output logic pcen,
						output logic [1:0]	pcsrc,
						output logic aluop
						output logic branch,
						output logic pcwrite);
						
						
	
				 
  
  
endmodule